ghjhjhujuhjhjhjhjhj