`default_nettype none
`timescale 1ns/1ns

module lsu(
    input wire clk,
    input wire reset,
    input wire enable,

    input reg [2:0] core_state,

     

);