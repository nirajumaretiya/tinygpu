`default_nettype none
`timescale 1ns/1ns

module controller #(
   parameter ADDR_BITS = 8,
   parameter DATA_BITS = 16,
   parameter NUM_CONSUMERS = 4,
   parameter NUM_CHANNELS= 1,
   parameter WRITE_ENABLE=1
)(
    input wire clk,
    input wire reset,
    
    input 
);

endmodule
